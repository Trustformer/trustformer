Require Import Koika.Frontend.
Require Import Koika.Std.
Require Koika.KoikaForm.Untyped.UntypedSemantics.
Require Import Koika.KoikaForm.SimpleVal.

Require Import Trustformer.v2_2.Syntax.
Require Import Trustformer.v2_2.Semantics.
Require Import Trustformer.v2_2.Synthesis.

Require Import Hammer.Plugin.Hammer.
Set Hammer GSMode 63.

(*
    An example specification and synthesis of a simple negator module.
    The hardware module has a single internal state register (32 bits) and supports two actions (nop, neg).
    Actions are triggered through a command register, where the first 1 bit indicates if the command is valid,
    and the remaining bits indicate the action to perform.

 *)

Section FunctionalSpecification.

    Definition sz := 32.
    Definition bits_false := Bits.of_nat sz 0.
    Definition bits_true := Bits.neg (bits_false).

    Inductive fs_action :=
    | fs_act_nop
    | fs_act_neg
    .

    Inductive fs_states :=
    | fs_st_val
    .

    Inductive fs_inputs :=
    .

    Inductive fs_outputs :=
    .

    Definition fs_states_size (x: fs_states) : nat :=
    match x with
    | fs_st_val => sz
    end.

    Definition fs_inputs_size (x: fs_inputs) : nat := 
    match x with
    end.

    Definition fs_outputs_size (x: fs_outputs) : nat := 
    match x with
    end.

    Definition fs_states_t := tf_states_type fs_states fs_states_size. 

    Definition fs_states_init (x: fs_states) : (fs_states_t x) :=
    match x with
    | fs_st_val => Bits.zero
    end.

    Definition fs_transitions
        (act: fs_action)
        :
        (tf_ops fs_states fs_inputs fs_outputs)
        :=
        match act with
        | fs_act_nop => tf_nop _ _ _ 
        | fs_act_neg => tf_neg _ _ _ fs_st_val
        end.

    Definition fs_step := tf_op_step_commit fs_states _ fs_inputs fs_outputs fs_states_size fs_inputs_size.
    
    Section Examples.

        Definition s_init := ContextEnv.(create) fs_states_init.
        Example s_example : ContextEnv.(getenv) s_init fs_st_val = bits_false.
        Proof. reflexivity. Qed.

        Definition s1_trans := fs_transitions fs_act_nop.
        Definition s1_state := fs_step s_init (fun _ => Bits.zero) s1_trans.
        Example s1_example : ContextEnv.(getenv) s1_state fs_st_val = bits_false.
        Proof. ssimpl. Qed.
        
        Definition s2_trans := fs_transitions fs_act_neg.
        Definition s2_state := fs_step s_init (fun _ => Bits.zero) s2_trans.
        Example s2_example : ContextEnv.(getenv) s2_state fs_st_val = bits_true.
        Proof. 
            cbn -[vect_to_list]. sauto.
        Qed.

    End Examples.

End FunctionalSpecification.


Section Synthesis.

    Definition tf_ctx : TFSynthContext := {|
        tf_spec_states := fs_states;
        tf_spec_states_fin := _; 
        tf_spec_states_size := fs_states_size;
        tf_spec_states_init := fs_states_init;

        tf_spec_inputs := fs_inputs;
        tf_spec_inputs_fin := _;
        tf_spec_inputs_size := fs_inputs_size;

        tf_spec_outputs := fs_outputs;
        tf_spec_outputs_fin := _;
        tf_spec_outputs_size := fs_outputs_size;

        tf_spec_action := fs_action;
        tf_spec_action_fin := _; 
        tf_spec_action_ops := fs_transitions
    |}.

    Definition R := Synthesis.R tf_ctx.

    Definition r := Synthesis.r tf_ctx.

    Definition Sigma := Synthesis.Sigma tf_ctx.

    Definition rules := Synthesis.rules tf_ctx.

    Definition system_schedule := Synthesis.system_schedule tf_ctx.
    
    Definition ext_fn_specs := Synthesis.ext_fn_specs tf_ctx.

    Instance ext_fn_names : Show (ext_fn_t tf_ctx) := Synthesis.ext_fn_names tf_ctx.

    Definition checked_rules := tc_rules R Sigma rules.

    Definition package :=
      {| ip_koika := {| koika_reg_types := R;
                        koika_reg_names := Synthesis.reg_names tf_ctx;
                        koika_reg_init := r;
                        koika_ext_fn_types := Sigma;
                        koika_rules := checked_rules;
                        koika_rule_names := Synthesis.rule_names tf_ctx;
                        koika_rule_external := (fun _ => false);
                        koika_scheduler := system_schedule;
                        koika_module_name := "V2_2Example_InternalNegator" |};

      ip_sim := {| sp_ext_fn_specs fn := {| efs_name := show fn; efs_method := false |};
                  sp_prelude := None |};

      ip_verilog := {| vp_ext_fn_specs := ext_fn_specs |} |}.
    

End Synthesis.

(* Extraction *)

Definition prog := Interop.Backends.register package.
Set Extraction Output Directory "build".
Extraction "V2_2Example_InternalNegator.ml" prog.

